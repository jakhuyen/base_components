module seg_display (
    input i_clk,
    input i_rst,
    input i_digit
);

    always @ (posedge i_rst, posedge i_clk) begin


    end

    
endmodule